// JWT - the namespace for this library/module
module jwt

// Imports: use `crypto.hmac` and `crypto.sha*` for signing the tokens
import crypto.hmac
import crypto.sha256
import crypto.sha512

// Functions
// Each of these functions generates an HMAC signature using either SHA 224, 
// 256, 384 or 512. The functions require base64 encoded headers, base64 
// encoded claims and a secret key to sign the headers and claims with. They 
// return the signature of the encoded headers and claims as a byte array

// Sign the headers and claims with HMAC-SHA224
fn hmac224(
	encoded_headers string,
	encoded_claims string,
	secret_key string
) []byte {
	return hmac.new(
		// The secret key
		secret_key.bytes(),
		// The content to sign
		(encoded_headers + '.' + encoded_claims).bytes(),
		// The function used to generate the checksum (here, SHA 224)
		sha256.sum224,
		// The size of a single block generated by the checksum function
		sha256.block_size
	)
}

// Sign the headers and claims with HMAC-SHA256
fn hmac256(
	encoded_headers string,
	encoded_claims string,
	secret_key string
) []byte {
	return hmac.new(
		// The secret key
		secret_key.bytes(),
		// The content to sign
		(encoded_headers + '.' + encoded_claims).bytes(),
		// The function used to generate the checksum (here, SHA 256)
		sha256.sum256,
		// The size of a single block generated by the checksum functions
		sha256.block_size
	)
}

// Sign the headers and claims with HMAC-SHA384
fn hmac384(
	encoded_headers string,
	encoded_claims string,
	secret_key string
) []byte {
	return hmac.new(
		// The secret key
		secret_key.bytes(),
		// The content to sign
		(encoded_headers + '.' + encoded_claims).bytes(),
		// The function used to generate the checksum (here, SHA 384)
		sha512.sum384,
		// The size of a single block generated by the checksum functions
		sha512.block_size
	)
}

// Sign the headers and claims with HMAC-SHA512
fn hmac512(
	encoded_headers string,
	encoded_claims string,
	secret_key string
) []byte {
	return hmac.new(
		// The secret key
		secret_key.bytes(),
		// The content to sign
		(encoded_headers + '.' + encoded_claims).bytes(),
		// The function used to generate the checksum (here, SHA 512/384)
		sha512.sum512_256,
		// The size of a single block generated by the checksum functions
		sha512.block_size
	)
}
